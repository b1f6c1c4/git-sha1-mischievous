`define METRIC 8 // $clog2(160+1)
`define BLOCKS 1
